magic
tech sky130A
timestamp 1739626261
<< nwell >>
rect 20 -145 195 0
rect 20 -155 180 -145
<< nmos >>
rect 95 -245 110 -195
<< pmos >>
rect 95 -135 110 -85
<< ndiff >>
rect 60 -205 95 -195
rect 60 -235 65 -205
rect 85 -235 95 -205
rect 60 -245 95 -235
rect 110 -205 145 -195
rect 110 -235 120 -205
rect 140 -235 145 -205
rect 110 -245 145 -235
<< pdiff >>
rect 60 -95 95 -85
rect 60 -125 65 -95
rect 85 -125 95 -95
rect 60 -135 95 -125
rect 110 -95 145 -85
rect 110 -125 120 -95
rect 140 -125 145 -95
rect 110 -135 145 -125
<< ndiffc >>
rect 65 -235 85 -205
rect 120 -235 140 -205
<< pdiffc >>
rect 65 -125 85 -95
rect 120 -125 140 -95
<< psubdiff >>
rect 60 -355 80 -330
rect 125 -355 145 -330
<< nsubdiff >>
rect 60 -45 80 -20
rect 120 -45 145 -20
<< psubdiffcont >>
rect 80 -355 125 -330
<< nsubdiffcont >>
rect 80 -45 120 -20
<< poly >>
rect 95 -85 110 -70
rect -5 -155 40 -150
rect 95 -155 110 -135
rect 160 -155 205 -150
rect -5 -175 5 -155
rect 25 -175 110 -155
rect 140 -175 175 -155
rect 195 -175 205 -155
rect -5 -180 40 -175
rect 95 -195 110 -175
rect 160 -180 205 -175
rect 95 -265 110 -245
<< polycont >>
rect 5 -175 25 -155
rect 175 -175 195 -155
<< locali >>
rect 60 -50 80 -20
rect 120 -45 145 -20
rect 60 -85 85 -50
rect 60 -95 90 -85
rect 60 -125 65 -95
rect 85 -125 90 -95
rect 60 -135 90 -125
rect 115 -95 145 -85
rect 115 -125 120 -95
rect 140 -125 145 -95
rect 115 -135 145 -125
rect -5 -155 40 -150
rect 120 -155 140 -135
rect 160 -155 205 -150
rect -5 -175 5 -155
rect 25 -175 90 -155
rect 120 -175 175 -155
rect 195 -175 205 -155
rect -5 -180 40 -175
rect 120 -195 140 -175
rect 160 -180 205 -175
rect 60 -205 90 -195
rect 60 -235 65 -205
rect 85 -235 90 -205
rect 60 -245 90 -235
rect 115 -205 145 -195
rect 115 -235 120 -205
rect 140 -235 145 -205
rect 115 -245 145 -235
rect 65 -330 90 -245
rect 60 -355 80 -330
rect 125 -355 145 -330
<< viali >>
rect 80 -20 120 -15
rect 80 -45 120 -20
rect 80 -50 120 -45
rect 5 -175 25 -155
rect 175 -175 195 -155
rect 80 -355 125 -330
<< metal1 >>
rect -10 -15 215 -10
rect -10 -50 80 -15
rect 120 -50 215 -15
rect -10 -55 215 -50
rect -5 -150 40 -145
rect -55 -155 40 -150
rect 160 -150 205 -145
rect 160 -155 255 -150
rect -55 -175 5 -155
rect 25 -175 95 -155
rect 120 -175 175 -155
rect 195 -175 255 -155
rect -55 -180 40 -175
rect -5 -185 40 -180
rect 160 -180 255 -175
rect 160 -185 205 -180
rect -10 -330 215 -325
rect -10 -355 80 -330
rect 125 -355 215 -330
rect -10 -360 215 -355
<< labels >>
rlabel metal1 180 -35 180 -35 1 vdd
rlabel metal1 180 -345 180 -345 1 vss
rlabel metal1 -35 -165 -35 -165 1 in
rlabel metal1 230 -165 230 -165 1 out
<< end >>
