** sch_path: /home/subramanian/VLSI projects/CMOS/inv_vtc.sch
**.subckt inv_vtc vdd vout vin gnd
*.ipin vin
*.ipin vdd
*.opin vout
*.ipin gnd
XM1 vout vin gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((1 + 1)/2) * 1 / 1 * 0.29' as='int((1 + 2)/2) * 1 / 1 * 0.29'
+ pd='2*int((1 + 1)/2) * (1 / 1 + 0.29)' ps='2*int((1 + 2)/2) * (1 / 1 + 0.29)' nrd='0.29 / 1 ' nrs='0.29 / 1 ' sa=0 sb=0 sd=0 mult=1
+ m=1
XM2 vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((1 + 1)/2) * 2 / 1 * 0.29' as='int((1 + 2)/2) * 2 / 1 * 0.29'
+ pd='2*int((1 + 1)/2) * (2 / 1 + 0.29)' ps='2*int((1 + 2)/2) * (2 / 1 + 0.29)' nrd='0.29 / 2 ' nrs='0.29 / 2 ' sa=0 sb=0 sd=0 mult=1
+ m=1
**.ends
.end
