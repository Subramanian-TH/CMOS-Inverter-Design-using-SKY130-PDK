magic
tech sky130A
timestamp 1765119862
<< nwell >>
rect -100 -150 200 260
<< nmos >>
rect 45 -355 60 -245
<< pmos >>
rect 45 -100 60 100
<< ndiff >>
rect -5 -255 45 -245
rect -5 -345 5 -255
rect 30 -345 45 -255
rect -5 -355 45 -345
rect 60 -255 110 -245
rect 60 -345 75 -255
rect 100 -345 110 -255
rect 60 -355 110 -345
<< pdiff >>
rect -5 90 45 100
rect -5 -90 5 90
rect 30 -90 45 90
rect -5 -100 45 -90
rect 60 90 110 100
rect 60 -90 75 90
rect 100 -90 110 90
rect 60 -100 110 -90
<< ndiffc >>
rect 5 -345 30 -255
rect 75 -345 100 -255
<< pdiffc >>
rect 5 -90 30 90
rect 75 -90 100 90
<< psubdiff >>
rect -10 -400 115 -385
rect -10 -425 5 -400
rect 100 -425 115 -400
rect -10 -440 115 -425
<< nsubdiff >>
rect -45 225 130 240
rect -45 205 -30 225
rect 115 205 130 225
rect -45 190 130 205
<< psubdiffcont >>
rect 5 -425 100 -400
<< nsubdiffcont >>
rect -30 205 115 225
<< poly >>
rect 45 100 60 160
rect 45 -150 60 -100
rect -15 -160 60 -150
rect -15 -185 -5 -160
rect 25 -185 60 -160
rect -15 -195 60 -185
rect 120 -160 170 -150
rect 120 -185 130 -160
rect 160 -185 170 -160
rect 120 -195 170 -185
rect 45 -245 60 -195
rect 45 -370 60 -355
<< polycont >>
rect -5 -185 25 -160
rect 130 -185 160 -160
<< locali >>
rect -45 225 130 240
rect -45 205 -30 225
rect 115 205 130 225
rect -45 190 130 205
rect 5 100 30 190
rect -5 90 40 100
rect -5 -90 5 90
rect 30 -90 40 90
rect -5 -100 40 -90
rect 65 90 110 100
rect 65 -90 75 90
rect 100 -90 110 90
rect 65 -100 110 -90
rect 75 -150 100 -100
rect -15 -160 35 -150
rect -15 -185 -5 -160
rect 25 -185 35 -160
rect -15 -195 35 -185
rect 75 -160 170 -150
rect 75 -185 130 -160
rect 160 -185 170 -160
rect 75 -195 170 -185
rect 75 -245 100 -195
rect -5 -255 40 -245
rect -5 -345 5 -255
rect 30 -345 40 -255
rect -5 -355 40 -345
rect 65 -255 110 -245
rect 65 -345 75 -255
rect 100 -345 110 -255
rect 65 -355 110 -345
rect 5 -390 30 -355
rect -5 -400 110 -390
rect -5 -425 5 -400
rect 100 -425 110 -400
rect -5 -435 110 -425
<< viali >>
rect 30 205 70 225
rect -5 -185 25 -160
rect 130 -185 160 -160
rect 35 -425 70 -400
<< metal1 >>
rect -165 225 250 240
rect -165 205 30 225
rect 70 205 250 225
rect -165 190 250 205
rect -130 -160 35 -150
rect -130 -185 -5 -160
rect 25 -185 35 -160
rect -130 -195 35 -185
rect 75 -160 235 -150
rect 75 -185 130 -160
rect 160 -185 235 -160
rect 75 -195 235 -185
rect -75 -400 185 -385
rect -75 -425 35 -400
rect 70 -425 185 -400
rect -75 -440 185 -425
<< labels >>
rlabel metal1 215 210 220 215 1 vdd
rlabel metal1 160 -410 165 -405 1 vss
rlabel metal1 195 -180 200 -175 1 out
rlabel metal1 -115 -185 -110 -180 1 in
<< end >>
